
module clk_div(clk,rst,div_clk);
    input clk,rst;
    output div_clk;
    reg div_clk;

    always @(posedge clk or negedge rst)
    begin
        if(!rst)
        begin
            div_clk <= 1'b0;
        end
        else
        begin
            div_clk = ~div_clk;
        end
    end
endmodule

module VGA_control(clk, rst, but_R, but_G, but_B, out_R, out_G, out_B,Hsync,Vsync);
    input clk, rst, but_R, but_G, but_B;
    output reg[3:0] out_R, out_G, out_B;
    output reg Hsync, Vsync;
    reg [9:0]counter_x, counter_y;
    reg [3:0]tmp_r,tmp_g,tmp_b;
    // counter and sync generation
    always @(posedge clk) // horizontal counter
    begin
        if(counter_x < 10'd799)
        begin
            counter_x <= counter_x + 10'd1; // horizontal counter (including off-screen horizontal 160 pixels) total of 800 pixels counter_x = 0~799
        end
        else
        begin
            counter_x <= 10'd0;
        end
    end // always

    always @ (posedge clk)  // vertical counter
    begin 
        if(counter_x == 10'd799)  // only counts up 1 count after horizontal finishes 800 counts
        begin
            if(counter_y < 10'd525) // vertical counter (including off-screen vertical 45 pixels) total of 525 pixels
            begin 
                counter_y <= counter_y + 10'd1;
            end
            else 
            begin
                counter_y <= 10'd0;
            end							 
        end  
    end  
    // end counter and sync generation  

    always @(posedge clk or negedge rst) 
    begin
        if(!rst)
        begin
            out_R <= 4'd0;
            out_G <= 4'd0;
            out_B <= 4'd0;
        end
        else 
        begin
            Hsync <= (counter_x >= 10'd0 && counter_x < 10'd96) ? 1'b0:1'b1;  // hsync low for 96 counts                                                 
            Vsync <= (counter_y >= 10'd0 && counter_y < 10'd2) ? 1'b0:1'b1;   // vsync low for 2 counts
            if(counter_x>=10'd96 && counter_x<=10'd144)
            begin               out_R <= 4'd0;
                out_G <= 4'd0;
                out_B <= 4'd0;
            end
            else
            begin
                out_R <= tmp_r;
                out_G <= tmp_g;
                out_B <= tmp_b;
            end
        end
	end
        
    
    always @(posedge but_R ) begin
        tmp_r <= tmp_r + 4'd1;
    end      
    always @(posedge but_G ) begin
        tmp_g <= tmp_g + 4'd1;
    end      
    always @(posedge but_B ) begin
        tmp_b <= tmp_b + 4'd1;
	end

    // assign Hsync = (counter_x >= 10'd0 && counter_x < 10'd96) ? 1'b0:1'b1;  // hsync low for 96 counts                                                 
    // assign Vsync = (counter_y >= 10'd0 && counter_y < 10'd2) ? 1'b0:1'b1;   // vsync low for 2 counts
endmodule


module VGA_display(clk, rst, num1,num2,num3,num4,num5,num6,num7,num8,num9,num10, enb, out_R, out_G, out_B,Hsync,Vsync);
    input clk, rst,enb;
    input [3:0]num1,num2,num3,num4,num5,num6,num7,num8,num9,num10;
    output reg[3:0] out_R, out_G, out_B;
    output reg Hsync, Vsync;
    reg [9:0]counter_x, counter_y;
    reg [3:0]tmp_r,tmp_g,tmp_b;
    // reg [31:0]old_num;
    // reg [3:0]num1;
    // reg [3:0]num2;
    // reg [3:0]num3;
    // reg [3:0]num4;
    // reg [3:0]num5;
    // reg [3:0]num6;
    // reg [3:0]num7;
    // reg [3:0]num8;
    // reg [3:0]num9;
    // reg [3:0]num10;

    // reg [3:0]tmp_num1;
    // reg [3:0]tmp_num2;
    // reg [3:0]tmp_num3;
    // reg [3:0]tmp_num4;
    // reg [3:0]tmp_num5;
    // reg [3:0]tmp_num6;
    // reg [3:0]tmp_num7;
    // reg [3:0]tmp_num8;
    // reg [3:0]tmp_num9;
    // reg [3:0]tmp_num10;
    // reg [5:0]i;
    // reg [71:0]shift_reg;  
    localparam [2499:0] zero = {
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000011000000000000000000000000,
			50'b00000000000000000000111111111110000000000000000000,
			50'b00000000000000000011111111111111100000000000000000,
			50'b00000000000000000111111111111111110000000000000000,
			50'b00000000000000001111111111111111111000000000000000,
			50'b00000000000000011111111111111111111100000000000000,
			50'b00000000000000111111111111111111111100000000000000,
			50'b00000000000000111111111000001111111110000000000000,
			50'b00000000000001111111110000000111111110000000000000,
			50'b00000000000001111111100000000011111111000000000000,
			50'b00000000000001111111000000000011111111000000000000,
			50'b00000000000011111111000000000001111111000000000000,
			50'b00000000000011111111000000000001111111000000000000,
			50'b00000000000011111111000000000001111111100000000000,
			50'b00000000000011111110000000000001111111100000000000,
			50'b00000000000011111110000000000001111111100000000000,
			50'b00000000000011111110000000000001111111100000000000,
			50'b00000000000011111110000000000001111111100000000000,
			50'b00000000000111111110000000000001111111100000000000,
			50'b00000000000111111110000000000001111111100000000000,
			50'b00000000000111111110000000000001111111100000000000,
			50'b00000000000111111110000000000001111111100000000000,
			50'b00000000000011111110000000000001111111100000000000,
			50'b00000000000011111110000000000001111111100000000000,
			50'b00000000000011111110000000000001111111100000000000,
			50'b00000000000011111110000000000001111111100000000000,
			50'b00000000000011111110000000000001111111100000000000,
			50'b00000000000011111111000000000001111111000000000000,
			50'b00000000000011111111000000000001111111000000000000,
			50'b00000000000001111111000000000011111111000000000000,
			50'b00000000000001111111100000000011111111000000000000,
			50'b00000000000001111111100000000111111110000000000000,
			50'b00000000000000111111110000001111111110000000000000,
			50'b00000000000000111111111111111111111100000000000000,
			50'b00000000000000011111111111111111111100000000000000,
			50'b00000000000000001111111111111111111000000000000000,
			50'b00000000000000000111111111111111110000000000000000,
			50'b00000000000000000011111111111111100000000000000000,
			50'b00000000000000000001111111111110000000000000000000,
			50'b00000000000000000000000111110000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000

    };

    localparam [2499:0] one = {
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000111111111111111111111111100000000000000,
			50'b00000000000111111111111111111111111100000000000000,
			50'b00000000000111111111111111111111111100000000000000,
			50'b00000000000111111111111111111111111100000000000000,
			50'b00000000000111111111111111111111111100000000000000,
			50'b00000000000000000001111111111000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111110000000000000000000000,
			50'b00000000000000000001111111111111111111100000000000,
			50'b00000000000000000001111111111111111111100000000000,
			50'b00000000000000000001111111111111111111100000000000,
			50'b00000000000000000001111111111111111110000000000000,
			50'b00000000000000000001111111111111111000000000000000,
			50'b00000000000000000001111111111110000000000000000000,
			50'b00000000000000000001111111100000000000000000000000,
			50'b00000000000000000001111100000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000
    };

    localparam [2499:0] two = {
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000001111111111111111111111111111000000000,
			50'b00000000000001111111111111111111111111111000000000,
			50'b00000000000001111111111111111111111111110000000000,
			50'b00000000000001111111111111111111111111110000000000,
			50'b00000000000001111111111111111111111111110000000000,
			50'b00000000000001111111111111111111111111110000000000,
			50'b00000000000000000000000000000011111111110000000000,
			50'b00000000000000000000000000000011111111100000000000,
			50'b00000000000000000000000000000111111111100000000000,
			50'b00000000000000000000000000001111111111000000000000,
			50'b00000000000000000000000000111111111110000000000000,
			50'b00000000000000000000000001111111111100000000000000,
			50'b00000000000000000000000111111111111000000000000000,
			50'b00000000000000000000001111111111110000000000000000,
			50'b00000000000000000000111111111111100000000000000000,
			50'b00000000000000000001111111111110000000000000000000,
			50'b00000000000000000111111111111100000000000000000000,
			50'b00000000000000001111111111110000000000000000000000,
			50'b00000000000000011111111111100000000000000000000000,
			50'b00000000000000011111111111000000000000000000000000,
			50'b00000000000000111111111100000000000000000000000000,
			50'b00000000000001111111111000000000000000000000000000,
			50'b00000000000001111111110000000000000000000000000000,
			50'b00000000000001111111110000000000000000000000000000,
			50'b00000000000001111111100000000000000000000000000000,
			50'b00000000000011111111100000000000111111110000000000,
			50'b00000000000011111111100000000000111111110000000000,
			50'b00000000000011111111100000000000111111110000000000,
			50'b00000000000011111111100000000000111111110000000000,
			50'b00000000000001111111100000000001111111100000000000,
			50'b00000000000001111111110000000001111111100000000000,
			50'b00000000000001111111111000000111111111100000000000,
			50'b00000000000000111111111111111111111111000000000000,
			50'b00000000000000111111111111111111111111000000000000,
			50'b00000000000000011111111111111111111110000000000000,
			50'b00000000000000001111111111111111111100000000000000,
			50'b00000000000000000111111111111111111000000000000000,
			50'b00000000000000000001111111111111100000000000000000,
			50'b00000000000000000000001111111100000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000

    };

    localparam [2499:0] three = {
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000111111100000000000000000000,
			50'b00000000000000000001111111111111100000000000000000,
			50'b00000000000000000011111111111111111000000000000000,
			50'b00000000000000001111111111111111111100000000000000,
			50'b00000000000000011111111111111111111110000000000000,
			50'b00000000000000111111111111111111111111000000000000,
			50'b00000000000000111111111100000111111111100000000000,
			50'b00000000000001111111110000000011111111100000000000,
			50'b00000000000001111111110000000001111111110000000000,
			50'b00000000000011111111100000000000111111110000000000,
			50'b00000000000011111111100000000000111111110000000000,
			50'b00000000000011111111100000000000010000000000000000,
			50'b00000000000011111111000000000000000000000000000000,
			50'b00000000000011111111100000000000000000000000000000,
			50'b00000000000011111111100000000000000000000000000000,
			50'b00000000000001111111100000000000000000000000000000,
			50'b00000000000001111111110000000000000000000000000000,
			50'b00000000000000111111111000000000000000000000000000,
			50'b00000000000000011111111111111100000000000000000000,
			50'b00000000000000001111111111111100000000000000000000,
			50'b00000000000000000011111111111000000000000000000000,
			50'b00000000000000000001111111111000000000000000000000,
			50'b00000000000000000111111111111000000000000000000000,
			50'b00000000000000001111111111111000000000000000000000,
			50'b00000000000000011111111100000000000000000000000000,
			50'b00000000000000011111111000000000000000000000000000,
			50'b00000000000000111111111000000000000000000000000000,
			50'b00000000000000111111110000000000000000000000000000,
			50'b00000000000000111111110000000000111111100000000000,
			50'b00000000000000111111110000000000111111100000000000,
			50'b00000000000000111111111000000001111111100000000000,
			50'b00000000000000111111111100000011111111100000000000,
			50'b00000000000000011111111111011111111111000000000000,
			50'b00000000000000001111111111111111111111000000000000,
			50'b00000000000000001111111111111111111110000000000000,
			50'b00000000000000000111111111111111111100000000000000,
			50'b00000000000000000001111111111111111000000000000000,
			50'b00000000000000000000011111111111000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000

    };

    localparam [2499:0] four = {
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000111111000000000000000000000000000,
			50'b00000000000000000111111100000000000000000000000000,
			50'b00000000000000000111111100000000000000000000000000,
			50'b00000000000000000111111100000000000000000000000000,
			50'b00000000000000000111111100000000000000000000000000,
			50'b00000000000000000111111100000000000000000000000000,
			50'b00000000000000000111111100000000000000000000000000,
			50'b00000000000000000111111100000000000000000000000000,
			50'b00000000000010001111111100000000000000000000000000,
			50'b00000000000011111111111111111111111111111000000000,
			50'b00000000000011111111111111111111111111111000000000,
			50'b00000000000011111111111111111111111111111000000000,
			50'b00000000000011111111111111111111111111110000000000,
			50'b00000000000011111111111111111111111111110000000000,
			50'b00000000000011111111111111111111111111110000000000,
			50'b00000000000000000111111100000000011111110000000000,
			50'b00000000000000000111111100000000011111110000000000,
			50'b00000000000000000111111100000000111111100000000000,
			50'b00000000000000000111111100000001111111000000000000,
			50'b00000000000000000111111100000011111110000000000000,
			50'b00000000000000000111111100000011111110000000000000,
			50'b00000000000000000111111100000111111100000000000000,
			50'b00000000000000000111111100001111111000000000000000,
			50'b00000000000000000111111100001111111000000000000000,
			50'b00000000000000000111111100011111110000000000000000,
			50'b00000000000000000111111100111111100000000000000000,
			50'b00000000000000000111111101111111000000000000000000,
			50'b00000000000000000111111101111111000000000000000000,
			50'b00000000000000000111111111111110000000000000000000,
			50'b00000000000000000111111111111100000000000000000000,
			50'b00000000000000000111111111111100000000000000000000,
			50'b00000000000000000111111111111000000000000000000000,
			50'b00000000000000000111111111110000000000000000000000,
			50'b00000000000000000111111111100000000000000000000000,
			50'b00000000000000000111111111100000000000000000000000,
			50'b00000000000000000111111111000000000000000000000000,
			50'b00000000000000000111111110000000000000000000000000,
			50'b00000000000000000111111110000000000000000000000000,
			50'b00000000000000000111111100000000000000000000000000,
			50'b00000000000000000111111000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000

    };

    localparam [2499:0]five = {
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000111111110000000000000000000,
			50'b00000000000000000000011111111111110000000000000000,
			50'b00000000000000000001111111111111111100000000000000,
			50'b00000000000000000111111111111111111110000000000000,
			50'b00000000000000001111111111111111111111000000000000,
			50'b00000000000000001111111111111111111111100000000000,
			50'b00000000000000011111111100000111111111100000000000,
			50'b00000000000000111111111000000001111111110000000000,
			50'b00000000000000111111110000000000111111110000000000,
			50'b00000000000000111111110000000000111111110000000000,
			50'b00000000000001111111100000000000011111110000000000,
			50'b00000000000001111111100000000000000000000000000000,
			50'b00000000000001111111100000000000000000000000000000,
			50'b00000000000001111111100000000000000000000000000000,
			50'b00000000000001111111100000000000000000000000000000,
			50'b00000000000001111111100000000000000000000000000000,
			50'b00000000000001111111100000000000000000000000000000,
			50'b00000000000001111111110000000000000000000000000000,
			50'b00000000000000111111111000000000111111100000000000,
			50'b00000000000000111111111100000001111111100000000000,
			50'b00000000000000011111111111111111111111100000000000,
			50'b00000000000000001111111111111111111111100000000000,
			50'b00000000000000001111111111111111111111100000000000,
			50'b00000000000000000011111111111111111111100000000000,
			50'b00000000000000000001111111111111111111000000000000,
			50'b00000000000000000000011111111101111111000000000000,
			50'b00000000000000000000000000000001111111000000000000,
			50'b00000000000000000000000000000011111111000000000000,
			50'b00000000000000000000000000000011111111000000000000,
			50'b00000000000000000000000000000011111110000000000000,
			50'b00000000000000000000000000000011111110000000000000,
			50'b00000000000000011111111111111111111110000000000000,
			50'b00000000000000011111111111111111111110000000000000,
			50'b00000000000000011111111111111111111100000000000000,
			50'b00000000000000011111111111111111111100000000000000,
			50'b00000000000000011111111111111111111100000000000000,
			50'b00000000000000011111111111111111111100000000000000,
			50'b00000000000000011111111111111111111100000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000

    };

    localparam [2499:0]six = {
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000111111111000000000000000000000,
			50'b00000000000000000111111111111111000000000000000000,
			50'b00000000000000011111111111111111110000000000000000,
			50'b00000000000000111111111111111111111000000000000000,
			50'b00000000000001111111111111111111111100000000000000,
			50'b00000000000011111111111111111111111110000000000000,
			50'b00000000000111111111110000111111111111000000000000,
			50'b00000000001111111111000000001111111111000000000000,
			50'b00000000001111111110000000000111111111100000000000,
			50'b00000000001111111110000000000011111111100000000000,
			50'b00000000001111111100000000000011111111110000000000,
			50'b00000000011111111100000000000011111111110000000000,
			50'b00000000011111111100000000000001111111110000000000,
			50'b00000000011111111100000000000001111111110000000000,
			50'b00000000011111111100000000000001111111111000000000,
			50'b00000000001111111100000000000011111111111000000000,
			50'b00000000001111111110000000000011111111111000000000,
			50'b00000000001111111110000000000011111111111000000000,
			50'b00000000000111111111000000001111111111111000000000,
			50'b00000000000111111111110000011111111111111000000000,
			50'b00000000000011111111111111111111111111111000000000,
			50'b00000000000001111111111111111111111111111000000000,
			50'b00000000000000111111111111111111111111111000000000,
			50'b00000000000000001111111111111101111111111000000000,
			50'b00000000000000000011111111100001111111110000000000,
			50'b00000000000000000000000000000001111111110000000000,
			50'b00000000000000000000000000000001111111110000000000,
			50'b00000000000000000000000000000001111111110000000000,
			50'b00000000000000000000000000000011111111100000000000,
			50'b00000000001111111110000000000011111111100000000000,
			50'b00000000001111111111000000000111111111100000000000,
			50'b00000000000111111111000000001111111111000000000000,
			50'b00000000000111111111111001111111111110000000000000,
			50'b00000000000011111111111111111111111110000000000000,
			50'b00000000000001111111111111111111111100000000000000,
			50'b00000000000000111111111111111111110000000000000000,
			50'b00000000000000011111111111111111100000000000000000,
			50'b00000000000000000111111111111100000000000000000000,
			50'b00000000000000000000011111100000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000

    };

    localparam [2499:0]seven ={
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000001111111111100000000000000,
			50'b00000000000000000000000001111111111100000000000000,
			50'b00000000000000000000000001111111111000000000000000,
			50'b00000000000000000000000011111111111000000000000000,
			50'b00000000000000000000000011111111111000000000000000,
			50'b00000000000000000000000011111111111000000000000000,
			50'b00000000000000000000000011111111111000000000000000,
			50'b00000000000000000000000011111111110000000000000000,
			50'b00000000000000000000000111111111110000000000000000,
			50'b00000000000000000000000111111111110000000000000000,
			50'b00000000000000000000000111111111100000000000000000,
			50'b00000000000000000000000111111111100000000000000000,
			50'b00000000000000000000001111111111100000000000000000,
			50'b00000000000000000000001111111111000000000000000000,
			50'b00000000000000000000011111111111000000000000000000,
			50'b00000000000000000000011111111110000000000000000000,
			50'b00000000000000000000111111111110000000000000000000,
			50'b00000000000000000000111111111100000000000000000000,
			50'b00000000000000000001111111111100000000000000000000,
			50'b00000000000000000001111111111000000000000000000000,
			50'b00000000000000000011111111111000000000000000000000,
			50'b00000000000000000011111111110000000000000000000000,
			50'b00000000000000000111111111100000000000000000000000,
			50'b00000000000000001111111111000000000000000000000000,
			50'b00000000000000001111111111000000000000000000000000,
			50'b00000000000000011111111110000000000000000000000000,
			50'b00000000000000111111111100000000000000000000000000,
			50'b00000000000001111111111000000000000000000000000000,
			50'b00000000000011111111111111111111111111111100000000,
			50'b00000000001111111111111111111111111111111100000000,
			50'b00000000001111111111111111111111111111111100000000,
			50'b00000000001111111111111111111111111111111100000000,
			50'b00000000001111111111111111111111111111111100000000,
			50'b00000000001111111111111111111111111111111100000000,
			50'b00000000001111111111111111111111111111111100000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000

    } ;

    localparam [2499:0]eight ={
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000011111111111111100000000000000000,
			50'b00000000000000011111111111111111111000000000000000,
			50'b00000000000001111111111111111111111110000000000000,
			50'b00000000000011111111111111111111111111000000000000,
			50'b00000000000111111111111111111111111111100000000000,
			50'b00000000000111111111111111111111111111110000000000,
			50'b00000000001111111111111100111111111111110000000000,
			50'b00000000001111111111110000001111111111111000000000,
			50'b00000000011111111111100000000111111111111000000000,
			50'b00000000011111111111100000000011111111111000000000,
			50'b00000000011111111111000000000011111111111000000000,
			50'b00000000011111111111000000000011111111111000000000,
			50'b00000000011111111111000000000011111111111000000000,
			50'b00000000011111111111000000000011111111111000000000,
			50'b00000000011111111111000000000011111111111000000000,
			50'b00000000011111111111100000000011111111111000000000,
			50'b00000000001111111111100000000111111111110000000000,
			50'b00000000000111111111110000001111111111110000000000,
			50'b00000000000111111111111111111111111111100000000000,
			50'b00000000000011111111111111111111111111000000000000,
			50'b00000000000001111111111111111111111110000000000000,
			50'b00000000000000011111111111111111111000000000000000,
			50'b00000000000000111111111111111111111100000000000000,
			50'b00000000000001111111111111111111111110000000000000,
			50'b00000000000011111111111111111111111111000000000000,
			50'b00000000000111111111111000011111111111100000000000,
			50'b00000000000111111111110000000111111111100000000000,
			50'b00000000000111111111100000000111111111110000000000,
			50'b00000000001111111111100000000011111111110000000000,
			50'b00000000001111111111100000000011111111110000000000,
			50'b00000000001111111111100000000011111111110000000000,
			50'b00000000001111111111100000000111111111110000000000,
			50'b00000000000111111111110000000111111111110000000000,
			50'b00000000000111111111111000011111111111100000000000,
			50'b00000000000111111111111111111111111111100000000000,
			50'b00000000000011111111111111111111111111000000000000,
			50'b00000000000001111111111111111111111110000000000000,
			50'b00000000000000111111111111111111111100000000000000,
			50'b00000000000000011111111111111111111000000000000000,
			50'b00000000000000000011111111111111100000000000000000,
			50'b00000000000000000000000111110000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000

    } ;

    localparam [2499:0]nine = {
        50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000001111111111111000000000000000000,
			50'b00000000000000000111111111111111111000000000000000,
			50'b00000000000000011111111111111111111100000000000000,
			50'b00000000000000011111111111111111111110000000000000,
			50'b00000000000000111111111111111111111111000000000000,
			50'b00000000000001111111111110011111111111000000000000,
			50'b00000000000001111111110000000111111111100000000000,
			50'b00000000000011111111110000000011111111100000000000,
			50'b00000000000011111111100000000011111111100000000000,
			50'b00000000000111111111100000000011111111100000000000,
			50'b00000000000111111111000000000000000000000000000000,
			50'b00000000000111111111000000000000000000000000000000,
			50'b00000000000111111111000000000000000000000000000000,
			50'b00000000000111111111000000000000000000000000000000,
			50'b00000000000111111111000011111111110000000000000000,
			50'b00000000000111111111001111111111111000000000000000,
			50'b00000000000111111111111111111111111110000000000000,
			50'b00000000000111111111111111111111111111000000000000,
			50'b00000000000111111111111111111111111111000000000000,
			50'b00000000000111111111111111111111111111100000000000,
			50'b00000000000111111111111100011111111111100000000000,
			50'b00000000000111111111110000000111111111100000000000,
			50'b00000000000111111111110000000011111111110000000000,
			50'b00000000000111111111100000000011111111110000000000,
			50'b00000000000111111111100000000011111111110000000000,
			50'b00000000000111111111100000000011111111110000000000,
			50'b00000000000111111111100000000011111111110000000000,
			50'b00000000000111111111100000000011111111110000000000,
			50'b00000000000111111111100000000011111111110000000000,
			50'b00000000000111111111100000000011111111110000000000,
			50'b00000000000111111111100000000011111111110000000000,
			50'b00000000000111111111100000000011111111110000000000,
			50'b00000000000111111111100000000011111111100000000000,
			50'b00000000000011111111110000000011111111100000000000,
			50'b00000000000011111111110000000111111111100000000000,
			50'b00000000000001111111111100011111111111000000000000,
			50'b00000000000001111111111111111111111111000000000000,
			50'b00000000000000111111111111111111111110000000000000,
			50'b00000000000000011111111111111111111100000000000000,
			50'b00000000000000001111111111111111111000000000000000,
			50'b00000000000000000001111111111111000000000000000000,
			50'b00000000000000000000001111110000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000,
			50'b00000000000000000000000000000000000000000000000000

    };

    // counter and sync generation
    always @(posedge clk) // horizontal counter
    begin
        if(counter_x < 10'd799)
        begin
            counter_x <= counter_x + 10'd1; // horizontal counter (including off-screen horizontal 160 pixels) total of 800 pixels counter_x = 0~799
        end
        else
        begin
            counter_x <= 10'd0;
        end
    end // always

    always @ (posedge clk)  // vertical counter
    begin 
        if(counter_x == 10'd799)  // only counts up 1 count after horizontal finishes 800 counts
        begin
            if(counter_y < 10'd525) // vertical counter (including off-screen vertical 45 pixels) total of 525 pixels
            begin 
                counter_y <= counter_y + 10'd1;
            end
            else 
            begin
                counter_y <= 10'd0;
            end							 
        end  
    end  
    // end counter and sync generation  
    //signal control
    always @(posedge clk or negedge rst) 
    begin
        if(!rst)
        begin
            out_R <= 4'd0;
            out_G <= 4'd0;
            out_B <= 4'd0;
        end
        else 
        begin
            Hsync <= (counter_x >= 10'd0 && counter_x < 10'd96) ? 1'b0:1'b1;  // hsync low for 96 counts                                                 
            Vsync <= (counter_y >= 10'd0 && counter_y < 10'd2) ? 1'b0:1'b1;   // vsync low for 2 counts
            if(counter_x>=10'd96 && counter_x<=10'd144)
            begin               
                out_R <= 4'd0;
                out_G <= 4'd0;
                out_B <= 4'd0;
            end
            else
            begin
                out_R <= tmp_r;
                out_G <= tmp_g;
                out_B <= tmp_b;
            end
        end
	end

    //bin 2 BCD
    // always @(posedge clk)
    //     begin
    //         //initialize bcd to zero.
    //         if(i == 6'd0 && (old_num != num))
    //         begin
    //             shift_reg <= 72'd0;
    //             old_num <= num;
    //             shift_reg[31:0] <= num;
    //             i <= i + 6'd1;
    //         end
    //         else if(i<6'd33 && i>6'd0)
    //         begin
    //             if(tmp_num10 >= 4'd5) tmp_num10 <= tmp_num10 + 4'd3;
    //             if(tmp_num9 >= 4'd5) tmp_num9 <= tmp_num9 + 4'd3;
    //             if(tmp_num8 >= 4'd5) tmp_num8 <= tmp_num8 + 4'd3;
    //             if(tmp_num7 >= 4'd5) tmp_num7 <= tmp_num7 + 4'd3;
    //             if(tmp_num6 >= 4'd5) tmp_num6 <= tmp_num6 + 4'd3;
    //             if(tmp_num5 >= 4'd5) tmp_num5 <= tmp_num5 + 4'd3;
    //             if(tmp_num4 >= 4'd5) tmp_num4 <= tmp_num4 + 4'd3;
    //             if(tmp_num3 >= 4'd5) tmp_num3 <= tmp_num3 + 4'd3;
    //             if(tmp_num2 >= 4'd5) tmp_num2 <= tmp_num2 + 4'd3;
    //             if(tmp_num1 >= 4'd5) tmp_num1 <= tmp_num1 + 4'd3;

    //             shift_reg [71:32] <= {tmp_num10,tmp_num9,tmp_num8,tmp_num7,tmp_num6,tmp_num5,tmp_num4,tmp_num3,tmp_num2,tmp_num1};
    //             shift_reg <= shift_reg << 1;
    //             tmp_num10 <= shift_reg[71:68];
    //             tmp_num9 <= shift_reg[67:64];
    //             tmp_num8 <= shift_reg[63:60];
    //             tmp_num7 <= shift_reg[59:56];
    //             tmp_num6 <= shift_reg[55:52];
    //             tmp_num5 <= shift_reg[51:48];
    //             tmp_num4 <= shift_reg[47:44];
    //             tmp_num3 <= shift_reg[43:40];
    //             tmp_num2 <= shift_reg[39:36];
    //             tmp_num1 <= shift_reg[35:32];
    //             i <= i + 6'd1;
    //         end
    //         else
    //         begin
    //             i <= 6'd0;
    //             num10 <= tmp_num10;
    //             num9 <= tmp_num9;
    //             num8 <= tmp_num8;
    //             num7 <= tmp_num7;
    //             num6 <= tmp_num6;
    //             num5 <= tmp_num5;
    //             num4 <= tmp_num4;
    //             num3 <= tmp_num3;
    //             num2 <= tmp_num2;
    //             num1 <= tmp_num1;
    //         end
    //     end
    // //function
    

    
    // pattern generate
        always @ (posedge clk)
        begin
            ////////////////////////////////////////////////////////////////////////////////////// SECTION 1
            if (counter_y < 50)//space to top
                begin              
                    tmp_r <= 4'h0;    // black
                    tmp_b <= 4'h0;
                    tmp_g <= 4'h0;
                end  
            ////////////////////////////////////////////////////////////////////////////////////// END SECTION 1
            
            ////////////////////////////////////////////////////////////////////////////////////// SECTION 2
            else if (counter_y >= 50 && counter_y < 55)
                begin 
                    if (counter_x >= 195 && counter_x < 705)
                        begin 
                            tmp_r <= 4'hF;    // white
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end  
                    else
                        begin 
                            tmp_r <= 4'h0;    // black
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end  
                    end 
            ////////////////////////////////////////////////////////////////////////////////////// END SECTION 2
            //display_num
            ////////////////////////////////////////////////////////////////////////////////////// SECTION 3
            else if (counter_y >= 55 && counter_y < 105)
                begin   
                    if (counter_x >= 195 && counter_x < 200)
                        begin 
                            tmp_r <= 4'hF;    // white
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end   
                    else if (counter_x >= 200 && counter_x < 250) //num10
                        if(enb)
                            begin
                                case(num10)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end 
                    else if (counter_x >= 250 && counter_x < 300) //num9
                        if(enb)
                            begin
                                case(num9)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[2499-(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 300 && counter_x < 350) //num8
                        if(enb)
                            begin
                                case(num8)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 350 && counter_x < 400) //num7
                        if(enb)
                            begin
                                case(num7)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 400 && counter_x < 450) //num6
                        if(enb)
                            begin
                                case(num6)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 450 && counter_x < 500) //num5
                        if(enb)
                            begin
                                case(num5)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 500 && counter_x < 550) //num4
                        if(enb)
                            begin
                                case(num4)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 550 && counter_x < 600) //num3
                        if(enb)
                            begin
                                case(num3)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 600 && counter_x < 650) //num2
                        if(enb)
                            begin
                                case(num2)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 650 && counter_x < 700) //num1
                        if(enb)
                            begin
                                case(num1)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 700 && counter_x < 705)
                        begin 
                            tmp_r <= 4'hF;    // white
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end 
                    else 
                        begin
                            tmp_r <= 4'h0;    // black
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end  // else if (counter_x >= 604)
                end  
            ////////////////////////////////////////////////////////////////////////////////////// END SECTION 3
            
            ////////////////////////////////////////////////////////////////////////////////////// SECTION 4
            else if (counter_y >= 105 && counter_y < 110)
                begin 
                    if (counter_x >= 195 && counter_x < 705)
                        begin 
                            tmp_r <= 4'hF;    // white
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end  
                    else
                        begin 
                            tmp_r <= 4'h0;    // black
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end  
                end 
				
				/*	  
				else 
					begin 
						tmp_r <= 4'h0;    // black
                  tmp_b <= 4'h0;
						tmp_g <= 4'h0;
					end
				*/
				else if (counter_y >= 110 && counter_y < 146)
                begin
                    tmp_r <= 4'h0;    // black
                    tmp_b <= 4'h0;
                    tmp_g <= 4'h0;
                end
            ///////////////////////////////////////////////////////////////////////////////////// 789 SECTION
            
				else if (counter_y >= 146 && counter_y < 151)
                begin
                    if ((counter_x >= 285 && counter_x < 335) || (counter_x >= 383 && counter_x <= 433) || (counter_x >= 481 && counter_x < 531 )
								|| (counter_x >= 579 && counter_x < 629))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else 
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            else if (counter_y >= 151 && counter_y < 201)
                begin
                    if((counter_x >= 280 && counter_x < 285) || (counter_x >= 335 && counter_x < 340) || (counter_x >=378 && counter_x < 383) || (counter_x >= 433 && counter_x < 438)
                        || (counter_x >= 476 && counter_x < 481) || (counter_x >= 531 && counter_x < 536) || (counter_x >= 574 && counter_x < 579) || (counter_x >= 629 && counter_x < 634))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            else if (counter_y >= 201 && counter_y < 206)
                begin
                    if ((counter_x >= 285 && counter_x < 335) || (counter_x >= 383 && counter_x <= 433) || (counter_x >= 481 && counter_x < 531 ) || (counter_x >= 579 && counter_x < 629 ))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else 
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            ///////////////////////////////////////////////////////////////////////////////////// 456 SECTION
            else if (counter_y >= 206 && counter_y < 230)
                begin
                    tmp_r <= 4'h0;    // black(0)
                    tmp_b <= 4'h0;
                    tmp_g <= 4'h0;
                end
            else if (counter_y >= 230 && counter_y < 235)
                begin
                    if ((counter_x >= 285 && counter_x < 335) || (counter_x >= 383 && counter_x <= 433) || (counter_x >= 481 && counter_x < 531 )
								|| (counter_x >= 579 && counter_x < 629))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else 
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            else if (counter_y >= 235 && counter_y < 285)
                begin
                    if((counter_x >= 280 && counter_x < 285) || (counter_x >= 335 && counter_x < 340) || (counter_x >=378 && counter_x < 383) || (counter_x >= 433 && counter_x < 438)
                        || (counter_x >= 476 && counter_x < 481) || (counter_x >= 531 && counter_x < 536) || (counter_x >= 574 && counter_x < 579) || (counter_x >= 629 && counter_x < 634))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            else if (counter_y >= 285 && counter_y < 290)
                begin
                   if ((counter_x >= 285 && counter_x < 335) || (counter_x >= 383 && counter_x <= 433) || (counter_x >= 481 && counter_x < 531 ) || (counter_x >= 579 && counter_x < 629 ))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else 
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            ////////////////////////////////////////////////////////////////////////////////////// 123 SECTION
            else if (counter_y >= 290 && counter_y < 314)
                begin
                    tmp_r <= 4'h0;    // black(0)
                    tmp_b <= 4'h0;
                    tmp_g <= 4'h0;
                end
            else if (counter_y >= 314 && counter_y < 319)
                begin
                     if ((counter_x >= 285 && counter_x < 335) || (counter_x >= 383 && counter_x <= 433) || (counter_x >= 481 && counter_x < 531 )
								|| (counter_x >= 579 && counter_x < 629))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else 
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            else if (counter_y >= 319 && counter_y < 369)
                begin
                    if((counter_x >= 280 && counter_x < 285) || (counter_x >= 335 && counter_x < 340) || (counter_x >=378 && counter_x < 383) || (counter_x >= 433 && counter_x < 438)
                        || (counter_x >= 476 && counter_x < 481) || (counter_x >= 531 && counter_x < 536) || (counter_x >= 574 && counter_x < 579) || (counter_x >= 629 && counter_x < 634))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            else if (counter_y >= 369 && counter_y < 374)
                begin
                    if ((counter_x >= 285 && counter_x < 335) || (counter_x >= 383 && counter_x <= 433) || (counter_x >= 481 && counter_x < 531 ) || (counter_x >= 579 && counter_x < 629 ))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else 
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            ////////////////////////////////////////////////////////////////////////////////////// 0 SECTION
            else if (counter_y >= 374 && counter_y < 398)
                begin
                    tmp_r <= 4'h0;    // black(0)
                    tmp_b <= 4'h0;
                    tmp_g <= 4'h0;
                end
            else if (counter_y >= 398 && counter_y < 403)
                begin
                     if ((counter_x >= 285 && counter_x < 335) || (counter_x >= 383 && counter_x <= 433) || (counter_x >= 481 && counter_x < 531 )
								|| (counter_x >= 579 && counter_x < 629))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else 
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            else if (counter_y >= 403 && counter_y < 453)
                begin
                   if((counter_x >= 280 && counter_x < 285) || (counter_x >= 335 && counter_x < 340) || (counter_x >=378 && counter_x < 383) || (counter_x >= 433 && counter_x < 438)
                        || (counter_x >= 476 && counter_x < 481) || (counter_x >= 531 && counter_x < 536) || (counter_x >= 574 && counter_x < 579) || (counter_x >= 629 && counter_x < 634))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            else if (counter_y >= 453 && counter_y < 458)
                begin
                    if ((counter_x >= 285 && counter_x < 335) || (counter_x >= 383 && counter_x <= 433) || (counter_x >= 481 && counter_x < 531 ) || (counter_x >= 579 && counter_x < 629 ))
                        begin
                            tmp_r <= 4'hF;    // white(1)
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end
                    else 
                        begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end
                end
            //////////////////////////////////////////////////////////////////////////////////////
            else
                begin
                            tmp_r <= 4'h0;    // black(0)
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                end
	 end  // always
						
endmodule

module input_num (clk,rst,but,num,enb);
    input clk,rst,but;
    output reg[31:0]num;
    output reg enb;
	 reg [31:0]tmp_num;
    always @(posedge clk or negedge rst ) begin
        if(!rst)
        begin
            enb <= 1'b0;
            num <= 32'b0;
        end 
        else
        begin
            enb <= 1'b1;
            num <= tmp_num;
        end
    end
    
	 always @(posedge but or negedge rst)
	 begin
		if(!rst)
		begin
			tmp_num <= 32'd0;
		end
		else
		begin
			tmp_num <= tmp_num + 32'd1;
		end
	 end
endmodule

module num2bcd(num,clk, output_num0, output_num1, output_num2, output_num3, output_num4, output_num5, output_num6, output_num7, output_num8, output_num9);
    input [31:0] num;
    input clk;
    output reg [3:0]output_num0;
    output reg [3:0]output_num1;
    output reg [3:0]output_num2;
    output reg [3:0]output_num3;
    output reg [3:0]output_num4;
    output reg [3:0]output_num5;
    output reg [3:0]output_num6;
    output reg [3:0]output_num7;
    output reg [3:0]output_num8;
    output reg [3:0]output_num9;

    reg [31:0] temp_num;
    reg [3:0]inter_num0;
    reg [3:0]inter_num1;
    reg [3:0]inter_num2;
    reg [3:0]inter_num3;
    reg [3:0]inter_num4;
    reg [3:0]inter_num5;
    reg [3:0]inter_num6;
    reg [3:0]inter_num7;
    reg [3:0]inter_num8;
    reg [3:0]inter_num9;
    reg[31:0]old_num;


    reg[8:0]state; // 0 (wait)+ 1~32(convert BCD)
    

    always @(posedge clk)
    begin
        if(state == 9'd0 && num != old_num)
        begin
            temp_num <= num;
            old_num <= num;
            state <= 9'd1;
            //  4'b1111 mean don't show number on display
            output_num0 <= 4'b1111;
            output_num1 <= 4'b1111;
            output_num2 <= 4'b1111;
            output_num3 <= 4'b1111;
            output_num4 <= 4'b1111;
            output_num5 <= 4'b1111;
            output_num6 <= 4'b1111;
            output_num7 <= 4'b1111;
            output_num8 <= 4'b1111;
            output_num9 <= 4'b1111;

            inter_num0 <= 4'b0000;
            inter_num1 <= 4'b0000;
            inter_num2 <= 4'b0000;
            inter_num3 <= 4'b0000;
            inter_num4 <= 4'b0000;
            inter_num5 <= 4'b0000;
            inter_num6 <= 4'b0000;
            inter_num7 <= 4'b0000;
            inter_num8 <= 4'b0000;
            inter_num9 <= 4'b0000;
        end

        else if(9'd1 <= state && state <= 9'd32)
        begin
            if(inter_num9 >=4'd5)
                inter_num9 = inter_num9 + 4'd3;
            if(inter_num8 >=4'd5)
                inter_num8 = inter_num8 + 4'd3;
            if(inter_num7 >=4'd5)
                inter_num7 = inter_num7 + 4'd3;
            if(inter_num6 >=4'd5)
                inter_num6 = inter_num6 + 4'd3;
            if(inter_num5 >=4'd5)
                inter_num5 = inter_num5 + 4'd3;
            if(inter_num4 >=4'd5)
                inter_num4 = inter_num4 + 4'd3;
            if(inter_num3 >=4'd5)
                inter_num3 = inter_num3 + 4'd3;
            if(inter_num2 >=4'd5)
                inter_num2 = inter_num2 + 4'd3;
            if(inter_num1 >=4'd5)
                inter_num1 = inter_num1 + 4'd3;
            if(inter_num0 >=4'd5)
                inter_num0 = inter_num0 + 4'd3;
            
            inter_num9 = inter_num9 << 1;
            inter_num9[0] = inter_num8[3];
            // inter_num9 = {inter_num9[2:0], inter_num8[3]};
            
            inter_num8 = inter_num8 << 1;
            inter_num8[0] = inter_num7[3];
            
            inter_num7 = inter_num7 << 1;
            inter_num7[0] = inter_num6[3];
            
            inter_num6 = inter_num6 << 1;
            inter_num6[0] = inter_num5[3];

            inter_num5 = inter_num5 << 1;
            inter_num5[0] = inter_num4[3];


            inter_num4 = inter_num4 << 1;
            inter_num4[0] = inter_num3[3];

            inter_num3 = inter_num3 << 1;
            inter_num3[0] = inter_num2[3];
            
            inter_num2 = inter_num2 << 1;
            inter_num2[0] = inter_num1[3];
            
            inter_num1 = inter_num1 << 1;
            inter_num1[0] = inter_num0[3];

            inter_num0 = inter_num0 << 1;
            inter_num0[0] = temp_num[31];

            temp_num = temp_num << 1; 
            state = state + 9'd1;
            
            if(state == 9'd33)
            begin
                state <= 9'd0;
                output_num0 <= inter_num0;
                output_num1 <= inter_num1;
                output_num2 <= inter_num2;
                output_num3 <= inter_num3;
                output_num4 <= inter_num4;
                output_num5 <= inter_num5;
                output_num6 <= inter_num6;
                output_num7 <= inter_num7;
                output_num8 <= inter_num8;
                output_num9 <= inter_num9;
            end
        end
    end
endmodule


module Freq_div(clk,clk_div);
	input clk;
	output reg clk_div;
	reg [24:0]counter;
	always@(posedge clk) begin
		if (counter == 25'd25000) begin // 1000Hz  (50M / (desire frequency))/2
			clk_div = ~clk_div;
			counter = counter +1;
		end
		else if (counter == 25'd50000) begin  //(50M / (desire frequency))
			clk_div = ~clk_div;
			counter = 0;
		end
		else
			counter <= counter +1;
	end
endmodule


module Freq_div2(clk,clk_div);
	input clk;
	output reg clk_div;
	reg [24:0]counter;
	always@(posedge clk) begin
		if (counter == 25'd2500000) begin // 1000Hz  (50M / (desire frequency))/2
			clk_div = ~clk_div;
			counter = counter +1;
		end
		else if (counter == 25'd5000000) begin  //(50M / (desire frequency))
			clk_div = ~clk_div;
			counter = 0;
		end
		else
			counter <= counter +1;
	end
endmodule


module Checkkeypad(clk_div,reset,keypadRow,keypadCol,keypadBuf);
	input clk_div;
	input reset;
	input [3:0]keypadCol;
	output reg[3:0]keypadRow;
	output reg [3:0] keypadBuf;
	always@(posedge clk_div or negedge reset) begin
		if (!reset)
		begin
			keypadRow <= 4'b1111;
			keypadBuf <= 0;
		end
		else begin
			case ({keypadRow,keypadCol})
				8'b1110_1110: keypadBuf <= 5'h7;
				8'b1110_1101: keypadBuf <= 5'h4;
				8'b1110_1011: keypadBuf <= 5'h1;
				8'b1110_0111: keypadBuf <= 5'h0;
				
				8'b1101_1110: keypadBuf <= 5'h8;
				8'b1101_1101: keypadBuf <= 5'h5;
				8'b1101_1011: keypadBuf <= 5'h2;
				8'b1101_0111: keypadBuf <= 5'ha;
				
				8'b1011_1110: keypadBuf <= 5'h9;
				8'b1011_1101: keypadBuf <= 5'h6;
				8'b1011_1011: keypadBuf <= 5'h3;
				8'b1011_0111: keypadBuf <= 5'hb;
				
				8'b0111_1110: keypadBuf <= 5'hc;
				8'b0111_1101: keypadBuf <= 5'hd;
				8'b0111_1011: keypadBuf <= 5'he;
				8'b0111_0111: keypadBuf <= 5'hf;
				default: keypadBuf <= keypadBuf;
				
			endcase
			case(keypadRow)
				4'b1110: keypadRow <= 4'b1101;
				4'b1101:	keypadRow <= 4'b1011;
				4'b1011:	keypadRow <= 4'b0111;
				4'b0111:	keypadRow <= 4'b1110;
				default: keypadRow <= 4'b1110;
			endcase
		end
	end
endmodule

module calculate(clk_div,reset,keypadBuf,keypadCol,out,enb);
   input clk_div;
	input reset;
	input[3:0] keypadBuf;
	input [3:0]keypadCol;
    reg[31:0] parameter1;
    reg[31:0] parameter2;
    output reg[31:0] out;
    reg[1:0] operand;
    reg flag,flag2;
	 reg[2:0]counter;
    output reg enb;

	 always@(posedge clk_div or negedge reset) begin
			if (!reset)
			begin
					flag2 <= 0;
			end
			else
			begin
					if(keypadCol != 4'hf)
					begin
							flag2 <= 1;
							counter <= 0;
					end
					
					else
					begin
					
							counter <= counter + 1;
							if(counter == 7)begin
									flag2 <= 0;
							end
					
					end
					
			end
	 end
	 always@(posedge flag2 or negedge reset) begin
			if (!reset)
			begin
			
					flag = 0;
					parameter1 <= 0;
					parameter2 <= 0;
					operand <= 0;
					out <= 0;
					enb <= 0;
			end
			else
			begin
				enb <= 1;
						case (keypadBuf)
							 5'ha:
							 begin
								  operand <= 0;
								  flag <= 1;
							 end
							 5'hb:
							 begin
								  operand <= 1;
								  flag <= 1;
							 end
							 5'hc:
							 begin
								  operand <= 2;
								  flag <= 1;
							 end
							 5'hd:
							 begin
								  operand <= 3;
								  flag <= 1;
							 end
							 5'he:
								  case(operand)
										0:
											 out <= parameter1 + parameter2;
										1:
											 out <= parameter1 - parameter2;
										2:
											 out <= parameter1 * parameter2;
										3:
											 out <= parameter1 / parameter2;
								  endcase
							 default:
								 begin
									if(flag == 0)begin
										parameter1 <= parameter1 *10 + keypadBuf;
										out <= parameter1 *10 + keypadBuf;
									end
									else
									begin
										parameter2 <= parameter2 *10 + keypadBuf;
										out <= parameter2;
									end
								end
								  
						endcase
				  
				
			end
	
	end
	
	 
endmodule



module VGA_output(clk,rst,but_R,but_G,but_B,out_R,out_G,out_B,Hsync,Vsync,keypadCol,keypadRow);

		
		input clk,rst,but_R,but_G,but_B;
		output [3:0] out_R,out_G,out_B;
		output Hsync, Vsync;
		wire div_clk,clk_div,clk_div2,enb;
		wire [31:0]num;
		wire [3:0]num1,num2,num3,num4,num5,num6,num7,num8,num9,num10;
		
		input [3:0]keypadCol;
		output [3:0]keypadRow;
		wire [4:0]keypadBuf;
		
		Freq_div u_Freq_div(.clk(clk),.clk_div(clk_div));
		//Freq_div2 u_Freq_div2(.clk(clk),.clk_div(clk_div2));
		clk_div u_clk_div(.clk(clk),.rst(rst),.div_clk(div_clk));
		
		Checkkeypad(.clk_div(clk_div),.reset(rst),.keypadRow(keypadRow),.keypadCol(keypadCol),.keypadBuf(keypadBuf));
		calculate(.clk_div(div_clk),.reset(rst),.keypadBuf(keypadBuf),.keypadCol(keypadCol),.out(num),.enb(enb));
		
		//input_num u_input_num(.clk(clk),.rst(rst),.but(but_B),.num(num),.enb(enb));
		
		
		num2bcd u_num2bcd(.num(num),.clk(clk), .output_num0(num1), .output_num1(num2), .output_num2(num3), .output_num3(num4), .output_num4(num5), .output_num5(num6), .output_num6(num7), .output_num7(num8), .output_num8(num9), .output_num9(num10));
		VGA_display u_VGA_display(.clk(div_clk), .rst(rst), .num1(num1),.num2(num2),.num3(num3),.num4(num4),.num5(num5),.num6(num6),.num7(num7),.num8(num8),.num9(num9),.num10(num10), .enb(enb), .out_R(out_R), .out_G(out_G), .out_B(out_B),.Hsync(Hsync),.Vsync(Vsync));
		
		
endmodule

