module clk_div(clk,rst,div_clk);
    input clk,rst;
    output div_clk;
    reg div_clk;

    always @(posedge clk or negedge rst)
    begin
        if(!rst)
        begin
            div_clk <= 1'b0;
        end
        else
        begin
            div_clk = ~div_clk;
        end
    end
endmodule

module VGA_control(clk, rst, but_R, but_G, but_B, out_R, out_G, out_B,Hsync,Vsync);
    input clk, rst, but_R, but_G, but_B;
    output reg[3:0] out_R, out_G, out_B;
    output reg Hsync, Vsync;
    reg [9:0]counter_x, counter_y;
    reg [3:0]tmp_r,tmp_g,tmp_b;
    // counter and sync generation
    always @(posedge clk) // horizontal counter
    begin
        if(counter_x < 10'd799)
        begin
            counter_x <= counter_x + 10'd1; // horizontal counter (including off-screen horizontal 160 pixels) total of 800 pixels counter_x = 0~799
        end
        else
        begin
            counter_x <= 10'd0;
        end
    end // always

    always @ (posedge clk)  // vertical counter
    begin 
        if(counter_x == 10'd799)  // only counts up 1 count after horizontal finishes 800 counts
        begin
            if(counter_y < 10'd525) // vertical counter (including off-screen vertical 45 pixels) total of 525 pixels
            begin 
                counter_y <= counter_y + 10'd1;
            end
            else 
            begin
                counter_y <= 10'd0;
            end							 
        end  
    end  
    // end counter and sync generation  

    always @(posedge clk or negedge rst) 
    begin
        if(!rst)
        begin
            out_R <= 4'd0;
            out_G <= 4'd0;
            out_B <= 4'd0;
        end
        else 
        begin
            Hsync <= (counter_x >= 10'd0 && counter_x < 10'd96) ? 1'b0:1'b1;  // hsync low for 96 counts                                                 
            Vsync <= (counter_y >= 10'd0 && counter_y < 10'd2) ? 1'b0:1'b1;   // vsync low for 2 counts
            if(counter_x>=10'd96 && counter_x<=10'd144)
            begin               out_R <= 4'd0;
                out_G <= 4'd0;
                out_B <= 4'd0;
            end
            else
            begin
                out_R <= tmp_r;
                out_G <= tmp_g;
                out_B <= tmp_b;
            end
        end
	end
        
    
    always @(posedge but_R ) begin
        tmp_r <= tmp_r + 4'd1;
    end      
    always @(posedge but_G ) begin
        tmp_g <= tmp_g + 4'd1;
    end      
    always @(posedge but_B ) begin
        tmp_b <= tmp_b + 4'd1;
	end

    // assign Hsync = (counter_x >= 10'd0 && counter_x < 10'd96) ? 1'b0:1'b1;  // hsync low for 96 counts                                                 
    // assign Vsync = (counter_y >= 10'd0 && counter_y < 10'd2) ? 1'b0:1'b1;   // vsync low for 2 counts
endmodule


module VGA_display(clk, rst, num, enb, out_R, out_G, out_B,Hsync,Vsync);
    input clk, rst,enb;
    input [31:0] num;
    output reg[3:0] out_R, out_G, out_B;
    output reg Hsync, Vsync;
    reg [9:0]counter_x, counter_y;
    reg [3:0]tmp_r,tmp_g,tmp_b;
    reg [31:0]old_num;
    reg [3:0]num1;
    reg [3:0]num2;
    reg [3:0]num3;
    reg [3:0]num4;
    reg [3:0]num5;
    reg [3:0]num6;
    reg [3:0]num7;
    reg [3:0]num8;
    reg [3:0]num9;
    reg [3:0]num10;

    reg [3:0]tmp_num1;
    reg [3:0]tmp_num2;
    reg [3:0]tmp_num3;
    reg [3:0]tmp_num4;
    reg [3:0]tmp_num5;
    reg [3:0]tmp_num6;
    reg [3:0]tmp_num7;
    reg [3:0]tmp_num8;
    reg [3:0]tmp_num9;
    reg [3:0]tmp_num10;
    reg [5:0]i;
    reg [71:0]shift_reg;  
    localparam [2499:0] zero = {
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000001111100000000000000000000000,
        50'b00000000000000000001111111111110000000000000000000,
        50'b00000000000000000111111111111111000000000000000000,
        50'b00000000000000001111111111111111100000000000000000,
        50'b00000000000000011111111111111111110000000000000000,
        50'b00000000000000111111111111111111111000000000000000,
        50'b00000000000000111111111111111111111100000000000000,
        50'b00000000000001111111110000001111111100000000000000,
        50'b00000000000001111111100000000111111110000000000000,
        50'b00000000000011111111000000000111111110000000000000,
        50'b00000000000011111111000000000011111110000000000000,
        50'b00000000000011111110000000000011111111000000000000,
        50'b00000000000011111110000000000011111111000000000000,
        50'b00000000000111111110000000000001111111000000000000,
        50'b00000000000111111110000000000001111111000000000000,
        50'b00000000000111111110000000000001111111000000000000,
        50'b00000000000111111110000000000001111111000000000000,
        50'b00000000000111111110000000000001111111000000000000,
        50'b00000000000111111110000000000001111111100000000000,
        50'b00000000000111111110000000000001111111100000000000,
        50'b00000000000111111110000000000001111111100000000000,
        50'b00000000000111111110000000000001111111100000000000,
        50'b00000000000111111110000000000001111111000000000000,
        50'b00000000000111111110000000000001111111000000000000,
        50'b00000000000111111110000000000001111111000000000000,
        50'b00000000000111111110000000000001111111000000000000,
        50'b00000000000111111110000000000011111111000000000000,
        50'b00000000000011111110000000000011111111000000000000,
        50'b00000000000011111110000000000011111111000000000000,
        50'b00000000000011111111000000000011111110000000000000,
        50'b00000000000011111111000000000111111110000000000000,
        50'b00000000000001111111100000001111111110000000000000,
        50'b00000000000001111111110000011111111100000000000000,
        50'b00000000000000111111111111111111111100000000000000,
        50'b00000000000000111111111111111111111000000000000000,
        50'b00000000000000011111111111111111110000000000000000,
        50'b00000000000000001111111111111111100000000000000000,
        50'b00000000000000000111111111111111000000000000000000,
        50'b00000000000000000001111111111100000000000000000000,
        50'b00000000000000000000000011000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000
    };

    localparam [2499:0] one = {
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000111111111111111111111111100000000000,
        50'b00000000000000111111111111111111111111100000000000,
        50'b00000000000000111111111111111111111111100000000000,
        50'b00000000000000111111111111111111111111100000000000,
        50'b00000000000000111111111111111111111111100000000000,
        50'b00000000000000000000011111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000000000000001111111110000000000000000000,
        50'b00000000000111111111111111111110000000000000000000,
        50'b00000000000111111111111111111110000000000000000000,
        50'b00000000000111111111111111111110000000000000000000,
        50'b00000000000001111111111111111110000000000000000000,
        50'b00000000000000011111111111111110000000000000000000,
        50'b00000000000000000001111111111110000000000000000000,
        50'b00000000000000000000000111111110000000000000000000,
        50'b00000000000000000000000000111110000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000
    };

    localparam [2499:0] two = {
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000011111111111111111111111111110000000000000,
        50'b00000000011111111111111111111111111110000000000000,
        50'b00000000001111111111111111111111111110000000000000,
        50'b00000000001111111111111111111111111110000000000000,
        50'b00000000001111111111111111111111111110000000000000,
        50'b00000000001111111111111111111111111110000000000000,
        50'b00000000001111111111000000000000000000000000000000,
        50'b00000000000111111111000000000000000000000000000000,
        50'b00000000000111111111100000000000000000000000000000,
        50'b00000000000011111111110000000000000000000000000000,
        50'b00000000000001111111111100000000000000000000000000,
        50'b00000000000000111111111110000000000000000000000000,
        50'b00000000000000011111111111100000000000000000000000,
        50'b00000000000000001111111111110000000000000000000000,
        50'b00000000000000000111111111111100000000000000000000,
        50'b00000000000000000001111111111110000000000000000000,
        50'b00000000000000000000111111111111100000000000000000,
        50'b00000000000000000000001111111111110000000000000000,
        50'b00000000000000000000000111111111111000000000000000,
        50'b00000000000000000000000011111111111000000000000000,
        50'b00000000000000000000000000111111111100000000000000,
        50'b00000000000000000000000000011111111110000000000000,
        50'b00000000000000000000000000001111111110000000000000,
        50'b00000000000000000000000000001111111110000000000000,
        50'b00000000000000000000000000000111111110000000000000,
        50'b00000000001111111100000000000111111111000000000000,
        50'b00000000001111111100000000000111111111000000000000,
        50'b00000000001111111100000000000111111111000000000000,
        50'b00000000001111111100000000000111111111000000000000,
        50'b00000000000111111110000000000111111110000000000000,
        50'b00000000000111111110000000001111111110000000000000,
        50'b00000000000111111111100000011111111110000000000000,
        50'b00000000000011111111111111111111111100000000000000,
        50'b00000000000011111111111111111111111100000000000000,
        50'b00000000000001111111111111111111111000000000000000,
        50'b00000000000000111111111111111111110000000000000000,
        50'b00000000000000011111111111111111100000000000000000,
        50'b00000000000000000111111111111110000000000000000000,
        50'b00000000000000000000111111110000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000  
    };

    localparam [2499:0] three = {
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000111111100000000000000000000000,
        50'b00000000000000000111111111111110000000000000000000,
        50'b00000000000000011111111111111111000000000000000000,
        50'b00000000000000111111111111111111110000000000000000,
        50'b00000000000001111111111111111111111000000000000000,
        50'b00000000000011111111111111111111111100000000000000,
        50'b00000000000111111111100000111111111100000000000000,
        50'b00000000000111111111000000001111111110000000000000,
        50'b00000000001111111110000000001111111110000000000000,
        50'b00000000001111111100000000000111111111000000000000,
        50'b00000000001111111100000000000111111111000000000000,
        50'b00000000000000001000000000000111111111000000000000,
        50'b00000000000000000000000000000011111111000000000000,
        50'b00000000000000000000000000000111111111000000000000,
        50'b00000000000000000000000000000111111111000000000000,
        50'b00000000000000000000000000000111111110000000000000,
        50'b00000000000000000000000000001111111110000000000000,
        50'b00000000000000000000000000011111111100000000000000,
        50'b00000000000000000000111111111111111000000000000000,
        50'b00000000000000000000111111111111110000000000000000,
        50'b00000000000000000000011111111111000000000000000000,
        50'b00000000000000000000011111111110000000000000000000,
        50'b00000000000000000000011111111111100000000000000000,
        50'b00000000000000000000011111111111110000000000000000,
        50'b00000000000000000000000000111111111000000000000000,
        50'b00000000000000000000000000011111111000000000000000,
        50'b00000000000000000000000000011111111100000000000000,
        50'b00000000000000000000000000001111111100000000000000,
        50'b00000000000111111100000000001111111100000000000000,
        50'b00000000000111111100000000001111111100000000000000,
        50'b00000000000111111110000000011111111100000000000000,
        50'b00000000000111111111000000111111111100000000000000,
        50'b00000000000011111111111011111111111000000000000000,
        50'b00000000000011111111111111111111110000000000000000,
        50'b00000000000001111111111111111111110000000000000000,
        50'b00000000000000111111111111111111100000000000000000,
        50'b00000000000000011111111111111110000000000000000000,
        50'b00000000000000000011111111111000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000
    };

    localparam [2499:0] four = {
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000011111100000000000000000,
        50'b00000000000000000000000000111111100000000000000000,
        50'b00000000000000000000000000111111100000000000000000,
        50'b00000000000000000000000000111111100000000000000000,
        50'b00000000000000000000000000111111100000000000000000,
        50'b00000000000000000000000000111111100000000000000000,
        50'b00000000000000000000000000111111100000000000000000,
        50'b00000000000000000000000000111111100000000000000000,
        50'b00000000000000000000000000111111110001000000000000,
        50'b00000000011111111111111111111111111111000000000000,
        50'b00000000011111111111111111111111111111000000000000,
        50'b00000000011111111111111111111111111111000000000000,
        50'b00000000001111111111111111111111111111000000000000,
        50'b00000000001111111111111111111111111111000000000000,
        50'b00000000001111111111111111111111111111000000000000,
        50'b00000000001111111000000000111111100000000000000000,
        50'b00000000001111111000000000111111100000000000000000,
        50'b00000000000111111100000000111111100000000000000000,
        50'b00000000000011111110000000111111100000000000000000,
        50'b00000000000001111111000000111111100000000000000000,
        50'b00000000000001111111000000111111100000000000000000,
        50'b00000000000000111111100000111111100000000000000000,
        50'b00000000000000011111110000111111100000000000000000,
        50'b00000000000000011111110000111111100000000000000000,
        50'b00000000000000001111111000111111100000000000000000,
        50'b00000000000000000111111100111111100000000000000000,
        50'b00000000000000000011111110111111100000000000000000,
        50'b00000000000000000011111110111111100000000000000000,
        50'b00000000000000000001111111111111100000000000000000,
        50'b00000000000000000000111111111111100000000000000000,
        50'b00000000000000000000111111111111100000000000000000,
        50'b00000000000000000000011111111111100000000000000000,
        50'b00000000000000000000001111111111100000000000000000,
        50'b00000000000000000000000111111111100000000000000000,
        50'b00000000000000000000000111111111100000000000000000,
        50'b00000000000000000000000011111111100000000000000000,
        50'b00000000000000000000000001111111100000000000000000,
        50'b00000000000000000000000001111111100000000000000000,
        50'b00000000000000000000000000111111100000000000000000,
        50'b00000000000000000000000000011111100000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000
    };

    localparam [2499:0]five = {
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000001111111100000000000000000000000,
        50'b00000000000000001111111111111000000000000000000000,
        50'b00000000000000111111111111111110000000000000000000,
        50'b00000000000001111111111111111111100000000000000000,
        50'b00000000000011111111111111111111110000000000000000,
        50'b00000000000111111111111111111111110000000000000000,
        50'b00000000000111111111100000111111111000000000000000,
        50'b00000000001111111110000000011111111100000000000000,
        50'b00000000001111111100000000001111111100000000000000,
        50'b00000000001111111100000000001111111100000000000000,
        50'b00000000001111111000000000000111111110000000000000,
        50'b00000000000000000000000000000111111110000000000000,
        50'b00000000000000000000000000000111111110000000000000,
        50'b00000000000000000000000000000111111110000000000000,
        50'b00000000000000000000000000000111111110000000000000,
        50'b00000000000000000000000000000111111110000000000000,
        50'b00000000000000000000000000000111111110000000000000,
        50'b00000000000000000000000000001111111110000000000000,
        50'b00000000000111111100000000011111111100000000000000,
        50'b00000000000111111110000000111111111100000000000000,
        50'b00000000000111111111111111111111111000000000000000,
        50'b00000000000111111111111111111111110000000000000000,
        50'b00000000000111111111111111111111110000000000000000,
        50'b00000000000111111111111111111111000000000000000000,
        50'b00000000000011111111111111111110000000000000000000,
        50'b00000000000011111110111111111000000000000000000000,
        50'b00000000000011111110000000000000000000000000000000,
        50'b00000000000011111111000000000000000000000000000000,
        50'b00000000000011111111000000000000000000000000000000,
        50'b00000000000001111111000000000000000000000000000000,
        50'b00000000000001111111000000000000000000000000000000,
        50'b00000000000001111111111111111111111000000000000000,
        50'b00000000000001111111111111111111111000000000000000,
        50'b00000000000000111111111111111111111000000000000000,
        50'b00000000000000111111111111111111111000000000000000,
        50'b00000000000000111111111111111111111000000000000000,
        50'b00000000000000111111111111111111111000000000000000,
        50'b00000000000000111111111111111111111000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000
    };

    localparam [2499:0]six = {
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000011111111100000000000000000000,
        50'b00000000000000000011111111111111100000000000000000,
        50'b00000000000000001111111111111111111000000000000000,
        50'b00000000000000011111111111111111111100000000000000,
        50'b00000000000000111111111111111111111110000000000000,
        50'b00000000000001111111111111111111111111000000000000,
        50'b00000000000011111111111100001111111111100000000000,
        50'b00000000000011111111110000000011111111110000000000,
        50'b00000000000111111111100000000001111111110000000000,
        50'b00000000000111111111000000000001111111110000000000,
        50'b00000000001111111111000000000000111111110000000000,
        50'b00000000001111111111000000000000111111111000000000,
        50'b00000000001111111110000000000000111111111000000000,
        50'b00000000001111111110000000000000111111111000000000,
        50'b00000000011111111110000000000000111111111000000000,
        50'b00000000011111111111000000000000111111110000000000,
        50'b00000000011111111111000000000001111111110000000000,
        50'b00000000011111111111000000000001111111110000000000,
        50'b00000000011111111111110000000011111111100000000000,
        50'b00000000011111111111111000001111111111100000000000,
        50'b00000000011111111111111111111111111111000000000000,
        50'b00000000011111111111111111111111111110000000000000,
        50'b00000000011111111111111111111111111100000000000000,
        50'b00000000011111111110111111111111110000000000000000,
        50'b00000000001111111110000111111111000000000000000000,
        50'b00000000001111111110000000000000000000000000000000,
        50'b00000000001111111110000000000000000000000000000000,
        50'b00000000001111111110000000000000000000000000000000,
        50'b00000000000111111111000000000000000000000000000000,
        50'b00000000000111111111000000000001111111110000000000,
        50'b00000000000111111111100000000011111111110000000000,
        50'b00000000000011111111110000000011111111100000000000,
        50'b00000000000001111111111110011111111111100000000000,
        50'b00000000000001111111111111111111111111000000000000,
        50'b00000000000000111111111111111111111110000000000000,
        50'b00000000000000001111111111111111111100000000000000,
        50'b00000000000000000111111111111111111000000000000000,
        50'b00000000000000000000111111111111100000000000000000,
        50'b00000000000000000000000111111000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000
    };

    localparam [2499:0]seven ={
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000111111111110000000000000000000000000,
        50'b00000000000000111111111110000000000000000000000000,
        50'b00000000000000011111111110000000000000000000000000,
        50'b00000000000000011111111111000000000000000000000000,
        50'b00000000000000011111111111000000000000000000000000,
        50'b00000000000000011111111111000000000000000000000000,
        50'b00000000000000011111111111000000000000000000000000,
        50'b00000000000000001111111111000000000000000000000000,
        50'b00000000000000001111111111100000000000000000000000,
        50'b00000000000000001111111111100000000000000000000000,
        50'b00000000000000000111111111100000000000000000000000,
        50'b00000000000000000111111111100000000000000000000000,
        50'b00000000000000000111111111110000000000000000000000,
        50'b00000000000000000011111111110000000000000000000000,
        50'b00000000000000000011111111111000000000000000000000,
        50'b00000000000000000001111111111000000000000000000000,
        50'b00000000000000000001111111111100000000000000000000,
        50'b00000000000000000000111111111100000000000000000000,
        50'b00000000000000000000111111111110000000000000000000,
        50'b00000000000000000000011111111110000000000000000000,
        50'b00000000000000000000011111111111000000000000000000,
        50'b00000000000000000000001111111111000000000000000000,
        50'b00000000000000000000000111111111100000000000000000,
        50'b00000000000000000000000011111111110000000000000000,
        50'b00000000000000000000000011111111110000000000000000,
        50'b00000000000000000000000001111111111000000000000000,
        50'b00000000000000000000000000111111111100000000000000,
        50'b00000000000000000000000000011111111110000000000000,
        50'b00000000111111111111111111111111111111000000000000,
        50'b00000000111111111111111111111111111111110000000000,
        50'b00000000111111111111111111111111111111110000000000,
        50'b00000000111111111111111111111111111111110000000000,
        50'b00000000111111111111111111111111111111110000000000,
        50'b00000000111111111111111111111111111111110000000000,
        50'b00000000111111111111111111111111111111110000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000
    } ;

    localparam [2499:0]eight ={
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000111111111111111000000000000000000,
        50'b00000000000000011111111111111111111000000000000000,
        50'b00000000000001111111111111111111111110000000000000,
        50'b00000000000011111111111111111111111111000000000000,
        50'b00000000000111111111111111111111111111100000000000,
        50'b00000000001111111111111111111111111111100000000000,
        50'b00000000001111111111111100111111111111110000000000,
        50'b00000000011111111111110000001111111111110000000000,
        50'b00000000011111111111100000000111111111111000000000,
        50'b00000000011111111111000000000111111111111000000000,
        50'b00000000011111111111000000000011111111111000000000,
        50'b00000000011111111111000000000011111111111000000000,
        50'b00000000011111111111000000000011111111111000000000,
        50'b00000000011111111111000000000011111111111000000000,
        50'b00000000011111111111000000000011111111111000000000,
        50'b00000000011111111111000000000111111111111000000000,
        50'b00000000001111111111100000000111111111110000000000,
        50'b00000000001111111111110000001111111111100000000000,
        50'b00000000000111111111111111111111111111100000000000,
        50'b00000000000011111111111111111111111111000000000000,
        50'b00000000000001111111111111111111111110000000000000,
        50'b00000000000000011111111111111111111000000000000000,
        50'b00000000000000111111111111111111111100000000000000,
        50'b00000000000001111111111111111111111110000000000000,
        50'b00000000000011111111111111111111111111000000000000,
        50'b00000000000111111111111000011111111111100000000000,
        50'b00000000000111111111100000001111111111100000000000,
        50'b00000000001111111111100000000111111111100000000000,
        50'b00000000001111111111000000000111111111110000000000,
        50'b00000000001111111111000000000111111111110000000000,
        50'b00000000001111111111000000000111111111110000000000,
        50'b00000000001111111111100000000111111111110000000000,
        50'b00000000001111111111100000001111111111100000000000,
        50'b00000000000111111111111000011111111111100000000000,
        50'b00000000000111111111111111111111111111100000000000,
        50'b00000000000011111111111111111111111111000000000000,
        50'b00000000000001111111111111111111111110000000000000,
        50'b00000000000000111111111111111111111100000000000000,
        50'b00000000000000011111111111111111111000000000000000,
        50'b00000000000000000111111111111111000000000000000000,
        50'b00000000000000000000001111100000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000
    } ;

    localparam [2499:0]nine = {
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000011111111111110000000000000000000,
        50'b00000000000000011111111111111111100000000000000000,
        50'b00000000000000111111111111111111111000000000000000,
        50'b00000000000001111111111111111111111000000000000000,
        50'b00000000000011111111111111111111111100000000000000,
        50'b00000000000011111111111001111111111110000000000000,
        50'b00000000000111111111100000001111111110000000000000,
        50'b00000000000111111111000000001111111111000000000000,
        50'b00000000000111111111000000000111111111000000000000,
        50'b00000000000111111111000000000111111111100000000000,
        50'b00000000000000000000000000000011111111100000000000,
        50'b00000000000000000000000000000011111111100000000000,
        50'b00000000000000000000000000000011111111100000000000,
        50'b00000000000000000000000000000011111111100000000000,
        50'b00000000000000001111111111000011111111100000000000,
        50'b00000000000000011111111111110011111111100000000000,
        50'b00000000000001111111111111111111111111100000000000,
        50'b00000000000011111111111111111111111111100000000000,
        50'b00000000000011111111111111111111111111100000000000,
        50'b00000000000111111111111111111111111111100000000000,
        50'b00000000000111111111111000111111111111100000000000,
        50'b00000000000111111111100000001111111111100000000000,
        50'b00000000001111111111000000001111111111100000000000,
        50'b00000000001111111111000000000111111111100000000000,
        50'b00000000001111111111000000000111111111100000000000,
        50'b00000000001111111111000000000111111111100000000000,
        50'b00000000001111111111000000000111111111100000000000,
        50'b00000000001111111111000000000111111111100000000000,
        50'b00000000001111111111000000000111111111100000000000,
        50'b00000000001111111111000000000111111111100000000000,
        50'b00000000001111111111000000000111111111100000000000,
        50'b00000000001111111111000000000111111111100000000000,
        50'b00000000000111111111000000000111111111100000000000,
        50'b00000000000111111111000000001111111111000000000000,
        50'b00000000000111111111100000001111111111000000000000,
        50'b00000000000011111111111000111111111110000000000000,
        50'b00000000000011111111111111111111111110000000000000,
        50'b00000000000001111111111111111111111100000000000000,
        50'b00000000000000111111111111111111111000000000000000,
        50'b00000000000000011111111111111111110000000000000000,
        50'b00000000000000000011111111111110000000000000000000,
        50'b00000000000000000000001111110000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000,
        50'b00000000000000000000000000000000000000000000000000
    };

    // counter and sync generation
    always @(posedge clk) // horizontal counter
    begin
        if(counter_x < 10'd799)
        begin
            counter_x <= counter_x + 10'd1; // horizontal counter (including off-screen horizontal 160 pixels) total of 800 pixels counter_x = 0~799
        end
        else
        begin
            counter_x <= 10'd0;
        end
    end // always

    always @ (posedge clk)  // vertical counter
    begin 
        if(counter_x == 10'd799)  // only counts up 1 count after horizontal finishes 800 counts
        begin
            if(counter_y < 10'd525) // vertical counter (including off-screen vertical 45 pixels) total of 525 pixels
            begin 
                counter_y <= counter_y + 10'd1;
            end
            else 
            begin
                counter_y <= 10'd0;
            end							 
        end  
    end  
    // end counter and sync generation  
    //signal control
    always @(posedge clk or negedge rst) 
    begin
        if(!rst)
        begin
            out_R <= 4'd0;
            out_G <= 4'd0;
            out_B <= 4'd0;
        end
        else 
        begin
            Hsync <= (counter_x >= 10'd0 && counter_x < 10'd96) ? 1'b0:1'b1;  // hsync low for 96 counts                                                 
            Vsync <= (counter_y >= 10'd0 && counter_y < 10'd2) ? 1'b0:1'b1;   // vsync low for 2 counts
            if(counter_x>=10'd96 && counter_x<=10'd144)
            begin               
                out_R <= 4'd0;
                out_G <= 4'd0;
                out_B <= 4'd0;
            end
            else
            begin
                out_R <= tmp_r;
                out_G <= tmp_g;
                out_B <= tmp_b;
            end
        end
	end

    //bin 2 BCD
    always @(posedge clk)
        begin
            //initialize bcd to zero.
            if(i == 6'd0 && (old_num != num))
            begin
                shift_reg <= 72'd0;
                old_num <= num;
                shift_reg[31:0] <= num;
                i <= i + 6'd1;
            end
            else if(i<33 && i>0)
            begin
                if(tmp_num10 >= 5) tmp_num10 <= tmp_num10 + 4'd3;
                if(tmp_num9 >= 5) tmp_num9 <= tmp_num9 + 4'd3;
                if(tmp_num8 >= 5) tmp_num8 <= tmp_num8 + 4'd3;
                if(tmp_num7 >= 5) tmp_num7 <= tmp_num7 + 4'd3;
                if(tmp_num6 >= 5) tmp_num6 <= tmp_num6 + 4'd3;
                if(tmp_num5 >= 5) tmp_num5 <= tmp_num5 + 4'd3;
                if(tmp_num4 >= 5) tmp_num4 <= tmp_num4 + 4'd3;
                if(tmp_num3 >= 5) tmp_num3 <= tmp_num3 + 4'd3;
                if(tmp_num2 >= 5) tmp_num2 <= tmp_num2 + 4'd3;
                if(tmp_num1 >= 5) tmp_num1 <= tmp_num1 + 4'd3;

                shift_reg [71:32] <= {tmp_num10,tmp_num9,tmp_num8,tmp_num7,tmp_num6,tmp_num5,tmp_num4,tmp_num3,tmp_num2,tmp_num1};
                shift_reg <= shift_reg << 1;
                tmp_num10 <= shift_reg[71:68];
                tmp_num9 <= shift_reg[67:64];
                tmp_num8 <= shift_reg[63:60];
                tmp_num7 <= shift_reg[59:56];
                tmp_num6 <= shift_reg[55:52];
                tmp_num5 <= shift_reg[51:48];
                tmp_num4 <= shift_reg[47:44];
                tmp_num3 <= shift_reg[43:40];
                tmp_num2 <= shift_reg[39:36];
                tmp_num1 <= shift_reg[35:32];
                i <= i + 6'd1;
            end
            else
            begin
                i <= 6'd0;
                num10 <= tmp_num10;
                num9 <= tmp_num9;
                num8 <= tmp_num8;
                num7 <= tmp_num7;
                num6 <= tmp_num6;
                num5 <= tmp_num5;
                num4 <= tmp_num4;
                num3 <= tmp_num3;
                num2 <= tmp_num2;
                num1 <= tmp_num1;
            end
        end

    // pattern generate
        always @ (posedge clk)
        begin
            ////////////////////////////////////////////////////////////////////////////////////// SECTION 1
            if (counter_y < 50)//space to top
                begin              
                    tmp_r <= 4'h0;    // black
                    tmp_b <= 4'h0;
                    tmp_g <= 4'h0;
                end  
            ////////////////////////////////////////////////////////////////////////////////////// END SECTION 1
            
            ////////////////////////////////////////////////////////////////////////////////////// SECTION 2
            else if (counter_y >= 50 && counter_y < 55)
                begin 
                    if (counter_x >= 195 && counter_x < 705)
                        begin 
                            tmp_r <= 4'hF;    // white
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end  
                    else
                        begin 
                            tmp_r <= 4'h0;    // black
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end  
                    end 
            ////////////////////////////////////////////////////////////////////////////////////// END SECTION 2
            //display_num
            ////////////////////////////////////////////////////////////////////////////////////// SECTION 3
            else if (counter_y >= 55 && counter_y < 105)
                begin   
                    if (counter_x >= 195 && counter_x < 200)
                        begin 
                            tmp_r <= 4'hF;    // white
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end   
                    else if (counter_x >= 200 && counter_x < 250)
                        begin 
                            if(enb)
                            begin
                                tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit10
                                tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // black
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                        end 
                    else if (counter_x >= 250 && counter_x < 300)
                        begin 
                            tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                            tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                            tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                        end
                    else if (counter_x >= 300 && counter_x < 350)
                        begin 
                            tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                            tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                            tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                        end
                    else if (counter_x >= 350 && counter_x < 400)
                        begin 
                            tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                            tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                            tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                        end
                    else if (counter_x >= 400 && counter_x < 450)
                        begin 
                            tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                            tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                            tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                        end
                    else if (counter_x >= 450 && counter_x < 500)
                        begin 
                            tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                            tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                            tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                        end
                    else if (counter_x >= 500 && counter_x < 550)
                        begin 
                            tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                            tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                            tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                        end
                    else if (counter_x >= 550 && counter_x < 600)
                        begin 
                            tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                            tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                            tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                        end
                    else if (counter_x >= 600 && counter_x < 650)
                        begin 
                            tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                            tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                            tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                        end
                    else if (counter_x >= 650 && counter_x < 700)
                        if(enb)
                            begin
                                case(num1)
                                    4'd0:
                                    begin
                                        tmp_r <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit0
                                        tmp_b <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (zero[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd1:
                                    begin
                                        tmp_r <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit1
                                        tmp_b <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (one[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd2:
                                    begin
                                        tmp_r <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit2
                                        tmp_b <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (two[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd3:
                                    begin
                                        tmp_r <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit3
                                        tmp_b <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (three[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd4:
                                    begin
                                        tmp_r <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit4
                                        tmp_b <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (four[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd5:
                                    begin
                                        tmp_r <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit5
                                        tmp_b <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (five[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd6:
                                    begin
                                        tmp_r <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit6
                                        tmp_b <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (six[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd7:
                                    begin
                                        tmp_r <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit7
                                        tmp_b <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (seven[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd8:
                                    begin
                                        tmp_r <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit8
                                        tmp_b <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (eight[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                    4'd9:
                                    begin
                                        tmp_r <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;    // digit9
                                        tmp_b <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                        tmp_g <= (nine[(counter_y-55)*50+(counter_x-300)]) ? 4'hF:4'h0;
                                    end
                                endcase
                            end
                            else
                            begin
                                tmp_r <= 4'h0;    // blank
                                tmp_b <= 4'h0;
                                tmp_g <= 4'h0;
                            end
                    else if (counter_x >= 700 && counter_x < 705)
                        begin 
                            tmp_r <= 4'hF;    // white
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end 
                    else 
                        begin
                            tmp_r <= 4'h0;    // black
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end  // else if (counter_x >= 604)
                end  
            ////////////////////////////////////////////////////////////////////////////////////// END SECTION 3
            
            ////////////////////////////////////////////////////////////////////////////////////// SECTION 4
            else if (counter_y >= 105 && counter_y < 110)
                begin 
                    if (counter_x >= 195 && counter_x < 705)
                        begin 
                            tmp_r <= 4'hF;    // white
                            tmp_b <= 4'hF;
                            tmp_g <= 4'hF;
                        end  
                    else
                        begin 
                            tmp_r <= 4'h0;    // black
                            tmp_b <= 4'h0;
                            tmp_g <= 4'h0;
                        end  
                end 
						  
				else 
					begin 
						tmp_r <= 4'h0;    // black
                  tmp_b <= 4'h0;
						tmp_g <= 4'h0;
					end
	 end  // always
						
	// end pattern generate
    // assign Hsync = (counter_x >= 10'd0 && counter_x < 10'd96) ? 1'b0:1'b1;  // hsync low for 96 counts                                                 
    // assign Vsync = (counter_y >= 10'd0 && counter_y < 10'd2) ? 1'b0:1'b1;   // vsync low for 2 counts
endmodule

module input_num (clk,rst,but,num,enb);
    input clk,rst,but;
    output reg[31:0]num;
    output reg enb;
    always @(posedge clk or negedge rst or posedge but) begin
        if(!rst)
        begin
            enb <= 1'b0;
            num <= 32'b0;
        end 
        else
        begin
            enb <= 1'b1;
            if(but)
            begin
                num <= num + 32'd1;
            end
            else
            begin 
                num <= num;
            end
        end
    end    
endmodule

module VGA_output(clk,rst,but_R,but_G,but_B,out_R,out_G,out_B,Hsync,Vsync);
    input clk,rst,but_R,but_G,but_B;
    output [3:0] out_R,out_G,out_B;
    output Hsync, Vsync;
    wire div_clk,enb;
    wire [31:0]num;
    clk_div u_clk_div(.clk(clk),.rst(rst),.div_clk(div_clk));
    input_num u_input_num(.clk(clk),.rst(rst),.but(but_B),.num(num),.enb(enb));
    VGA_display u_VGA_display(.clk(div_clk), .rst(rst), .num(num), .enb(enb), .out_R(out_R), .out_G(out_G), .out_B(out_B),.Hsync(Hsync),.Vsync(Vsync));
endmodule

